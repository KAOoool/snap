module  transform_memory(
                     clk,
                     rst,
                 i_valid,
              i_transize,
                     
                     i_0,
                     i_1,
                     i_2,
                     i_3,
                     i_4,
                     i_5,
                     i_6,
                     i_7,
                     i_8,
                     i_9,
                     i_10,
                     i_11,
                     i_12,
                     i_13,
                     i_14,
                     i_15,
                     i_16,
                     i_17,
                     i_18,
                     i_19,
                     i_20,
                     i_21,
                     i_22,
                     i_23,
                     i_24,
                     i_25,
                     i_26,
                     i_27,
                     i_28,
                     i_29,
                     i_30,
                     i_31,
                     
                  o_valid,
                      o_0, 
                      o_1,
                      o_2,
                      o_3,
					  o_4, 
					  o_5,
					  o_6,
				   	  o_7,
					  o_8, 
					  o_9,
					 o_10,
					 o_11,
					 o_12,
					 o_13,
					 o_14,
				   o_15,
					 o_16,
					 o_17,
					 o_18,
					 o_19,
					 o_20,
					 o_21,
					 o_22,
					 o_23,
					 o_24,
					 o_25,
					 o_26,
					 o_27,
					 o_28,
				 	 o_29,
					 o_30,
					 o_31
);
                     
// ********************************************
//                                             
//    INPUT / OUTPUT DECLARATION                                               
//                                                                             
// ********************************************

input                         clk;
input                         rst;
input                     i_valid;
input signed [1:0]     i_transize;
input signed [15:0]           i_0;
input signed [15:0]           i_1;
input signed [15:0]           i_2;
input signed [15:0]           i_3;
input signed [15:0]           i_4;
input signed [15:0]           i_5;
input signed [15:0]           i_6;
input signed [15:0]           i_7;
input signed [15:0]           i_8;
input signed [15:0]           i_9;
input signed [15:0]           i_10;
input signed [15:0]           i_11;
input signed [15:0]           i_12;
input signed [15:0]           i_13;
input signed [15:0]           i_14;
input signed [15:0]           i_15;
input signed [15:0]           i_16;
input signed [15:0]           i_17;
input signed [15:0]           i_18;
input signed [15:0]           i_19;
input signed [15:0]           i_20;
input signed [15:0]           i_21;
input signed [15:0]           i_22;
input signed [15:0]           i_23;
input signed [15:0]           i_24;
input signed [15:0]           i_25;
input signed [15:0]           i_26;
input signed [15:0]           i_27;
input signed [15:0]           i_28;
input signed [15:0]           i_29;
input signed [15:0]           i_30;
input signed [15:0]           i_31;

output  reg                o_valid;
output signed [15:0]           o_0; 
output signed [15:0]           o_1;
output signed [15:0]           o_2;
output signed [15:0]           o_3;
output signed [15:0]           o_4; 
output signed [15:0]           o_5;
output signed [15:0]           o_6;
output signed [15:0]           o_7;
output signed [15:0]           o_8; 
output signed [15:0]           o_9;
output signed [15:0]           o_10;
output signed [15:0]           o_11;
output signed [15:0]           o_12; 
output signed [15:0]           o_13;
output signed [15:0]           o_14;
output signed [15:0]           o_15;
output signed [15:0]           o_16; 
output signed [15:0]           o_17;
output signed [15:0]           o_18;
output signed [15:0]           o_19;
output signed [15:0]           o_20; 
output signed [15:0]           o_21;
output signed [15:0]           o_22;
output signed [15:0]           o_23;
output signed [15:0]           o_24; 
output signed [15:0]           o_25;
output signed [15:0]           o_26;
output signed [15:0]           o_27;
output signed [15:0]           o_28; 
output signed [15:0]           o_29;
output signed [15:0]           o_30;
output signed [15:0]           o_31;


// ********************************************
//                                             
//    Wire DECLARATION                         
//                                             
// ********************************************
wire                              wen;
wire                           enable;
wire         [4:0]            counter;

wire         [4:0]            badd_0 ;
wire         [4:0]            badd_1 ;
wire         [4:0]            badd_2 ;
wire         [4:0]            badd_3 ;
wire         [4:0]            badd_4 ;
wire         [4:0]            badd_5 ;
wire         [4:0]            badd_6 ;
wire         [4:0]            badd_7 ;
wire         [4:0]            badd_8 ;
wire         [4:0]            badd_9 ;
wire         [4:0]            badd_10;
wire         [4:0]            badd_11;
wire         [4:0]            badd_12;
wire         [4:0]            badd_13;
wire         [4:0]            badd_14;
wire         [4:0]            badd_15;
wire         [4:0]            badd_16;
wire         [4:0]            badd_17;
wire         [4:0]            badd_18;
wire         [4:0]            badd_19;
wire         [4:0]            badd_20;
wire         [4:0]            badd_21;
wire         [4:0]            badd_22;
wire         [4:0]            badd_23;
wire         [4:0]            badd_24;
wire         [4:0]            badd_25;
wire         [4:0]            badd_26;
wire         [4:0]            badd_27;
wire         [4:0]            badd_28;
wire         [4:0]            badd_29;
wire         [4:0]            badd_30;
wire         [4:0]            badd_31;
wire         [4:0]             add_0 ;
wire         [4:0]             add_1 ;
wire         [4:0]             add_2 ;
wire         [4:0]             add_3 ;
wire         [4:0]             add_4 ;
wire         [4:0]             add_5 ;
wire         [4:0]             add_6 ;
wire         [4:0]             add_7 ;
wire         [4:0]             add_8 ;
wire         [4:0]             add_9 ;
wire         [4:0]             add_10;
wire         [4:0]             add_11;
wire         [4:0]             add_12;
wire         [4:0]             add_13;
wire         [4:0]             add_14;
wire         [4:0]             add_15;
wire         [4:0]             add_16;
wire         [4:0]             add_17;
wire         [4:0]             add_18;
wire         [4:0]             add_19;
wire         [4:0]             add_20;
wire         [4:0]             add_21;
wire         [4:0]             add_22;
wire         [4:0]             add_23;
wire         [4:0]             add_24;
wire         [4:0]             add_25;
wire         [4:0]             add_26;
wire         [4:0]             add_27;
wire         [4:0]             add_28;
wire         [4:0]             add_29;
wire         [4:0]             add_30;
wire         [4:0]             add_31;

wire signed  [15:0]           i_m_0 ;
wire signed  [15:0]           i_m_1 ;
wire signed  [15:0]           i_m_2 ;
wire signed  [15:0]           i_m_3 ;
wire signed  [15:0]           i_m_4 ;
wire signed  [15:0]           i_m_5 ;
wire signed  [15:0]           i_m_6 ;
wire signed  [15:0]           i_m_7 ;
wire signed  [15:0]           i_m_8 ;
wire signed  [15:0]           i_m_9 ;
wire signed  [15:0]           i_m_10;
wire signed  [15:0]           i_m_11;
wire signed  [15:0]           i_m_12;
wire signed  [15:0]           i_m_13;
wire signed  [15:0]           i_m_14;
wire signed  [15:0]           i_m_15;
wire signed  [15:0]           i_m_16;
wire signed  [15:0]           i_m_17;
wire signed  [15:0]           i_m_18;
wire signed  [15:0]           i_m_19;
wire signed  [15:0]           i_m_20;
wire signed  [15:0]           i_m_21;
wire signed  [15:0]           i_m_22;
wire signed  [15:0]           i_m_23;
wire signed  [15:0]           i_m_24;
wire signed  [15:0]           i_m_25;
wire signed  [15:0]           i_m_26;
wire signed  [15:0]           i_m_27;
wire signed  [15:0]           i_m_28;
wire signed  [15:0]           i_m_29;
wire signed  [15:0]           i_m_30;
wire signed  [15:0]           i_m_31;

wire signed  [15:0]           o_m_0 ;
wire signed  [15:0]           o_m_1 ;
wire signed  [15:0]           o_m_2 ;
wire signed  [15:0]           o_m_3 ;
wire signed  [15:0]           o_m_4 ;
wire signed  [15:0]           o_m_5 ;
wire signed  [15:0]           o_m_6 ;
wire signed  [15:0]           o_m_7 ;
wire signed  [15:0]           o_m_8 ;
wire signed  [15:0]           o_m_9 ;
wire signed  [15:0]           o_m_10;
wire signed  [15:0]           o_m_11;
wire signed  [15:0]           o_m_12;
wire signed  [15:0]           o_m_13;
wire signed  [15:0]           o_m_14;
wire signed  [15:0]           o_m_15;
wire signed  [15:0]           o_m_16;
wire signed  [15:0]           o_m_17;
wire signed  [15:0]           o_m_18;
wire signed  [15:0]           o_m_19;
wire signed  [15:0]           o_m_20;
wire signed  [15:0]           o_m_21;
wire signed  [15:0]           o_m_22;
wire signed  [15:0]           o_m_23;
wire signed  [15:0]           o_m_24;
wire signed  [15:0]           o_m_25;
wire signed  [15:0]           o_m_26;
wire signed  [15:0]           o_m_27;
wire signed  [15:0]           o_m_28;
wire signed  [15:0]           o_m_29;
wire signed  [15:0]           o_m_30;
wire signed  [15:0]           o_m_31;


wire signed  [15:0]           i_s_0 ;
wire signed  [15:0]           i_s_1 ;
wire signed  [15:0]           i_s_2 ;
wire signed  [15:0]           i_s_3 ;
wire signed  [15:0]           i_s_4 ;
wire signed  [15:0]           i_s_5 ;
wire signed  [15:0]           i_s_6 ;
wire signed  [15:0]           i_s_7 ;
wire signed  [15:0]           i_s_8 ;
wire signed  [15:0]           i_s_9 ;
wire signed  [15:0]           i_s_10;
wire signed  [15:0]           i_s_11;
wire signed  [15:0]           i_s_12;
wire signed  [15:0]           i_s_13;
wire signed  [15:0]           i_s_14;
wire signed  [15:0]           i_s_15;
wire signed  [15:0]           i_s_16;
wire signed  [15:0]           i_s_17;
wire signed  [15:0]           i_s_18;
wire signed  [15:0]           i_s_19;
wire signed  [15:0]           i_s_20;
wire signed  [15:0]           i_s_21;
wire signed  [15:0]           i_s_22;
wire signed  [15:0]           i_s_23;
wire signed  [15:0]           i_s_24;
wire signed  [15:0]           i_s_25;
wire signed  [15:0]           i_s_26;
wire signed  [15:0]           i_s_27;
wire signed  [15:0]           i_s_28;
wire signed  [15:0]           i_s_29;
wire signed  [15:0]           i_s_30;
wire signed  [15:0]           i_s_31;

wire signed  [15:0]           o_s_0 ;
wire signed  [15:0]           o_s_1 ;
wire signed  [15:0]           o_s_2 ;
wire signed  [15:0]           o_s_3 ;
wire signed  [15:0]           o_s_4 ;
wire signed  [15:0]           o_s_5 ;
wire signed  [15:0]           o_s_6 ;
wire signed  [15:0]           o_s_7 ;
wire signed  [15:0]           o_s_8 ;
wire signed  [15:0]           o_s_9 ;
wire signed  [15:0]           o_s_10;
wire signed  [15:0]           o_s_11;
wire signed  [15:0]           o_s_12;
wire signed  [15:0]           o_s_13;
wire signed  [15:0]           o_s_14;
wire signed  [15:0]           o_s_15;
wire signed  [15:0]           o_s_16;
wire signed  [15:0]           o_s_17;
wire signed  [15:0]           o_s_18;
wire signed  [15:0]           o_s_19;
wire signed  [15:0]           o_s_20;
wire signed  [15:0]           o_s_21;
wire signed  [15:0]           o_s_22;
wire signed  [15:0]           o_s_23;
wire signed  [15:0]           o_s_24;
wire signed  [15:0]           o_s_25;
wire signed  [15:0]           o_s_26;
wire signed  [15:0]           o_s_27;
wire signed  [15:0]           o_s_28;
wire signed  [15:0]           o_s_29;
wire signed  [15:0]           o_s_30;
wire signed  [15:0]           o_s_31;



// ********************************************
//                                             
//    Reg DECLARATION                         
//                                             
// ********************************************

reg                       o_chose;             
reg                         wen_0;
reg                         wen_1;
reg                      enable_0;

reg signed [15:0]           i_r_0;
reg signed [15:0]           i_r_1;
reg signed [15:0]           i_r_2;
reg signed [15:0]           i_r_3;
reg signed [15:0]           i_r_4;
reg signed [15:0]           i_r_5;
reg signed [15:0]           i_r_6;
reg signed [15:0]           i_r_7;
reg signed [15:0]           i_r_8;
reg signed [15:0]           i_r_9;
reg signed [15:0]           i_r_10;
reg signed [15:0]           i_r_11;
reg signed [15:0]           i_r_12;
reg signed [15:0]           i_r_13;
reg signed [15:0]           i_r_14;
reg signed [15:0]           i_r_15;
reg signed [15:0]           i_r_16;
reg signed [15:0]           i_r_17;
reg signed [15:0]           i_r_18;
reg signed [15:0]           i_r_19;
reg signed [15:0]           i_r_20;
reg signed [15:0]           i_r_21;
reg signed [15:0]           i_r_22;
reg signed [15:0]           i_r_23;
reg signed [15:0]           i_r_24;
reg signed [15:0]           i_r_25;
reg signed [15:0]           i_r_26;
reg signed [15:0]           i_r_27;
reg signed [15:0]           i_r_28;
reg signed [15:0]           i_r_29;
reg signed [15:0]           i_r_30;
reg signed [15:0]           i_r_31;

// ********************************************
//                                             
//    Combinational Logic                      
//                                             
// ********************************************

assign i_m_0 =wen_1?o_s_0 :i_0 ;
assign i_m_1 =wen_1?o_s_1 :i_1 ;
assign i_m_2 =wen_1?o_s_2 :i_2 ;
assign i_m_3 =wen_1?o_s_3 :i_3 ;
assign i_m_4 =wen_1?o_s_4 :i_4 ;
assign i_m_5 =wen_1?o_s_5 :i_5 ;
assign i_m_6 =wen_1?o_s_6 :i_6 ;
assign i_m_7 =wen_1?o_s_7 :i_7 ;
assign i_m_8 =wen_1?o_s_8 :i_8 ;
assign i_m_9 =wen_1?o_s_9 :i_9 ;
assign i_m_10=wen_1?o_s_10:i_10;
assign i_m_11=wen_1?o_s_11:i_11;
assign i_m_12=wen_1?o_s_12:i_12;
assign i_m_13=wen_1?o_s_13:i_13;
assign i_m_14=wen_1?o_s_14:i_14;
assign i_m_15=wen_1?o_s_15:i_15;
assign i_m_16=wen_1?o_s_16:i_16;
assign i_m_17=wen_1?o_s_17:i_17;
assign i_m_18=wen_1?o_s_18:i_18;
assign i_m_19=wen_1?o_s_19:i_19;
assign i_m_20=wen_1?o_s_20:i_20;
assign i_m_21=wen_1?o_s_21:i_21;
assign i_m_22=wen_1?o_s_22:i_22;
assign i_m_23=wen_1?o_s_23:i_23;
assign i_m_24=wen_1?o_s_24:i_24;
assign i_m_25=wen_1?o_s_25:i_25;
assign i_m_26=wen_1?o_s_26:i_26;
assign i_m_27=wen_1?o_s_27:i_27;
assign i_m_28=wen_1?o_s_28:i_28;
assign i_m_29=wen_1?o_s_29:i_29;
assign i_m_30=wen_1?o_s_30:i_30;
assign i_m_31=wen_1?o_s_31:i_31;

assign i_s_0 =wen_0?16'b0:o_m_0 ;
assign i_s_1 =wen_0?16'b0:o_m_1 ;
assign i_s_2 =wen_0?16'b0:o_m_2 ;
assign i_s_3 =wen_0?16'b0:o_m_3 ;
assign i_s_4 =wen_0?16'b0:o_m_4 ;
assign i_s_5 =wen_0?16'b0:o_m_5 ;
assign i_s_6 =wen_0?16'b0:o_m_6 ;
assign i_s_7 =wen_0?16'b0:o_m_7 ;
assign i_s_8 =wen_0?16'b0:o_m_8 ;
assign i_s_9 =wen_0?16'b0:o_m_9 ;
assign i_s_10=wen_0?16'b0:o_m_10;
assign i_s_11=wen_0?16'b0:o_m_11;
assign i_s_12=wen_0?16'b0:o_m_12;
assign i_s_13=wen_0?16'b0:o_m_13;
assign i_s_14=wen_0?16'b0:o_m_14;
assign i_s_15=wen_0?16'b0:o_m_15;
assign i_s_16=wen_0?16'b0:o_m_16;
assign i_s_17=wen_0?16'b0:o_m_17;
assign i_s_18=wen_0?16'b0:o_m_18;
assign i_s_19=wen_0?16'b0:o_m_19;
assign i_s_20=wen_0?16'b0:o_m_20;
assign i_s_21=wen_0?16'b0:o_m_21;
assign i_s_22=wen_0?16'b0:o_m_22;
assign i_s_23=wen_0?16'b0:o_m_23;
assign i_s_24=wen_0?16'b0:o_m_24;
assign i_s_25=wen_0?16'b0:o_m_25;
assign i_s_26=wen_0?16'b0:o_m_26;
assign i_s_27=wen_0?16'b0:o_m_27;
assign i_s_28=wen_0?16'b0:o_m_28;
assign i_s_29=wen_0?16'b0:o_m_29;
assign i_s_30=wen_0?16'b0:o_m_30;
assign i_s_31=wen_0?16'b0:o_m_31;

assign o_0  =o_chose?o_m_0: 16'b0;
assign o_1  =o_chose?o_m_1: 16'b0;
assign o_2  =o_chose?o_m_2: 16'b0;
assign o_3  =o_chose?o_m_3: 16'b0;
assign o_4  =o_chose?o_m_4: 16'b0;
assign o_5  =o_chose?o_m_5: 16'b0;
assign o_6  =o_chose?o_m_6: 16'b0;
assign o_7  =o_chose?o_m_7: 16'b0;
assign o_8  =o_chose?o_m_8: 16'b0;
assign o_9  =o_chose?o_m_9: 16'b0;
assign o_10 =o_chose?o_m_10:16'b0;
assign o_11 =o_chose?o_m_11:16'b0;
assign o_12 =o_chose?o_m_12:16'b0;
assign o_13 =o_chose?o_m_13:16'b0;
assign o_14 =o_chose?o_m_14:16'b0;
assign o_15 =o_chose?o_m_15:16'b0;
assign o_16 =o_chose?o_m_16:16'b0;
assign o_17 =o_chose?o_m_17:16'b0;
assign o_18 =o_chose?o_m_18:16'b0;
assign o_19 =o_chose?o_m_19:16'b0;
assign o_20 =o_chose?o_m_20:16'b0;
assign o_21 =o_chose?o_m_21:16'b0;
assign o_22 =o_chose?o_m_22:16'b0;
assign o_23 =o_chose?o_m_23:16'b0;
assign o_24 =o_chose?o_m_24:16'b0;
assign o_25 =o_chose?o_m_25:16'b0;
assign o_26 =o_chose?o_m_26:16'b0;
assign o_27 =o_chose?o_m_27:16'b0;
assign o_28 =o_chose?o_m_28:16'b0;
assign o_29 =o_chose?o_m_29:16'b0;
assign o_30 =o_chose?o_m_30:16'b0;
assign o_31 =o_chose?o_m_31:16'b0;

always@(*)
o_valid=o_chose;

// ********************************************
//                                             
//    Sequential  Logic                        
//                                             
// ********************************************

always@(posedge clk or negedge rst)
if(!rst)
o_chose<=1'b0;
else
  if(i_transize==2'b00)
    o_chose<=i_valid;
  else
    o_chose<=wen_1;

always@(posedge clk or negedge rst)
if(!rst)
 enable_0<=1'b0;
else
  enable_0<=enable;
   
always@(posedge clk or negedge rst)
if(!rst)
  wen_0<=1'b0;
else
  wen_0<=wen;

 always@(posedge clk or negedge rst)
if(!rst)
  wen_1<=1'b0;
else
  wen_1<=wen_0;
  
always@(posedge clk or negedge rst)
if(!rst)
begin
i_r_0<=16'b0;
i_r_1<=16'b0;
i_r_2<=16'b0; 
i_r_3<=16'b0; 
i_r_4<=16'b0; 
i_r_5<=16'b0; 
i_r_6<=16'b0; 
i_r_7<=16'b0; 
i_r_8<=16'b0; 
i_r_9<=16'b0; 
i_r_10<=16'b0; 
i_r_11<=16'b0; 
i_r_12<=16'b0; 
i_r_13<=16'b0; 
i_r_14<=16'b0; 
i_r_15<=16'b0; 
i_r_16<=16'b0; 
i_r_17<=16'b0; 
i_r_18<=16'b0; 
i_r_19<=16'b0; 
i_r_20<=16'b0; 
i_r_21<=16'b0; 
i_r_22<=16'b0; 
i_r_23<=16'b0; 
i_r_24<=16'b0; 
i_r_25<=16'b0; 
i_r_26<=16'b0; 
i_r_27<=16'b0; 
i_r_28<=16'b0; 
i_r_29<=16'b0; 
i_r_30<=16'b0; 
i_r_31<=16'b0; 
end
else
begin
 i_r_0 <= i_m_0 ;
 i_r_1 <= i_m_1 ;
 i_r_2 <= i_m_2 ;
 i_r_3 <= i_m_3 ;
 i_r_4 <= i_m_4 ;
 i_r_5 <= i_m_5 ;
 i_r_6 <= i_m_6 ;
 i_r_7 <= i_m_7 ;
 i_r_8 <= i_m_8 ;
 i_r_9 <= i_m_9 ;
 i_r_10<= i_m_10;
 i_r_11<= i_m_11;
 i_r_12<= i_m_12;
 i_r_13<= i_m_13;
 i_r_14<= i_m_14;
 i_r_15<= i_m_15;
 i_r_16<= i_m_16;
 i_r_17<= i_m_17;
 i_r_18<= i_m_18;
 i_r_19<= i_m_19;
 i_r_20<= i_m_20;
 i_r_21<= i_m_21;
 i_r_22<= i_m_22;
 i_r_23<= i_m_23;
 i_r_24<= i_m_24;
 i_r_25<= i_m_25;
 i_r_26<= i_m_26;
 i_r_27<= i_m_27;
 i_r_28<= i_m_28;
 i_r_29<= i_m_29;
 i_r_30<= i_m_30;
 i_r_31<= i_m_31;
 end
 
 
// ********************************************
//                                             
//    Sub Modules                              
//                                             
// ********************************************

ctrl_transmemory  ctrl_transmemory_0(
                    clk,
                    rst,
                i_valid,
             i_transize,
             
                    wen,
                 enable,
                counter
);

addr        add0_0(
              clk,
              rst,
           enable,
              wen,
          counter, 
       i_transize,
       
		      badd_0 ,
          badd_1 ,
          badd_2 ,
          badd_3 ,
          badd_4 ,
          badd_5 ,
          badd_6 ,
          badd_7 ,
          badd_8 ,
          badd_9 ,
          badd_10,
          badd_11,
          badd_12,
          badd_13,
          badd_14,
          badd_15,
          badd_16,
          badd_17,
          badd_18,
          badd_19,
          badd_20,
          badd_21,
          badd_22,
          badd_23,
          badd_24,
          badd_25,
          badd_26,
          badd_27,
          badd_28,
          badd_29,
          badd_30,
          badd_31,
           add_0 ,
           add_1 ,
           add_2 ,
           add_3 ,
           add_4 ,
           add_5 ,
           add_6 ,
           add_7 ,
           add_8 ,
           add_9 ,
           add_10,
           add_11,
           add_12,
           add_13,
           add_14,
           add_15,
           add_16,
           add_17,
           add_18,
           add_19,
           add_20,
           add_21,
           add_22,
           add_23,
           add_24,
           add_25,
           add_26,
           add_27,
           add_28,
           add_29,
           add_30,
           add_31
);
              
mux_32    mux_32_0(
              badd_0,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_0
);

mux_32    mux_32_1(
              badd_1,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_1
);

mux_32    mux_32_2(
              badd_2,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_2
);

mux_32    mux_32_3(
              badd_3,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_3
);

mux_32    mux_32_4(
              badd_4,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_4
);

mux_32    mux_32_5(
              badd_5,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_5
);

mux_32    mux_32_6(
              badd_6,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_6
);

mux_32    mux_32_7(
              badd_7,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_7
);

mux_32    mux_32_8(
              badd_8,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_8
);

mux_32    mux_32_9(
              badd_9,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_9
);

mux_32    mux_32_10(
             badd_10,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_10
);

mux_32    mux_32_11(
             badd_11,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_11
);

mux_32    mux_32_12(
             badd_12,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_12
);

mux_32    mux_32_13(
             badd_13,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
               o_m_13
);

mux_32    mux_32_14(
             badd_14,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_14
);

mux_32    mux_32_15(
             badd_15,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_15
);

mux_32    mux_32_16(
             badd_16,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_16
);

mux_32    mux_32_17(
             badd_17,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_17
);

mux_32    mux_32_18(
             badd_18,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_18
);

mux_32    mux_32_19(
             badd_19,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_19
);

mux_32    mux_32_20(
             badd_20,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_20
);

mux_32    mux_32_21(
             badd_21,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_21
);

mux_32    mux_32_22(
             badd_22,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_22
);

mux_32    mux_32_23(
             badd_23,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_23
);

mux_32    mux_32_24(
             badd_24,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_24
);

mux_32    mux_32_25(
             badd_25,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_25
);

mux_32    mux_32_26(
             badd_26,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_26
);

mux_32    mux_32_27(
             badd_27,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_27
);

mux_32    mux_32_28(
             badd_28,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_28
);

mux_32    mux_32_29(
             badd_29,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_29
);

mux_32    mux_32_30(
             badd_30,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_30
);

mux_32    mux_32_31(
             badd_31,
              i_r_0 ,
              i_r_1 ,
              i_r_2 ,
              i_r_3 ,
              i_r_4 ,
              i_r_5 ,
              i_r_6 ,
              i_r_7 ,
              i_r_8 ,
              i_r_9 ,
              i_r_10,
              i_r_11,
              i_r_12,
              i_r_13,
              i_r_14,
              i_r_15,
              i_r_16,
              i_r_17,
              i_r_18,
              i_r_19,
              i_r_20,
              i_r_21,
              i_r_22,
              i_r_23,
              i_r_24,
              i_r_25,
              i_r_26,
              i_r_27,
              i_r_28,
              i_r_29,
              i_r_30,
              i_r_31,
          
              o_m_31
);

tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_0(.data_o(o_s_0),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_0),.data_i(i_s_0),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_1(.data_o(o_s_1),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_1),.data_i(i_s_1),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_2(.data_o(o_s_2),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_2),.data_i(i_s_2),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_3(.data_o(o_s_3),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_3),.data_i(i_s_3),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_4(.data_o(o_s_4),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_4),.data_i(i_s_4),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_5(.data_o(o_s_5),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_5),.data_i(i_s_5),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_6(.data_o(o_s_6),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_6),.data_i(i_s_6),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_7(.data_o(o_s_7),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_7),.data_i(i_s_7),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_8(.data_o(o_s_8),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_8),.data_i(i_s_8),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_9(.data_o(o_s_9),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_9),.data_i(i_s_9),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_10(.data_o(o_s_10),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_10),.data_i(i_s_10),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_11(.data_o(o_s_11),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_11),.data_i(i_s_11),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_12(.data_o(o_s_12),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_12),.data_i(i_s_12),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_13(.data_o(o_s_13),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_13),.data_i(i_s_13),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_14(.data_o(o_s_14),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_14),.data_i(i_s_14),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_15(.data_o(o_s_15),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_15),.data_i(i_s_15),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_16(.data_o(o_s_16),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_16),.data_i(i_s_16),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_17(.data_o(o_s_17),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_17),.data_i(i_s_17),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_18(.data_o(o_s_18),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_18),.data_i(i_s_18),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_19(.data_o(o_s_19),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_19),.data_i(i_s_19),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_20(.data_o(o_s_20),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_20),.data_i(i_s_20),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_21(.data_o(o_s_21),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_21),.data_i(i_s_21),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_22(.data_o(o_s_22),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_22),.data_i(i_s_22),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_23(.data_o(o_s_23),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_23),.data_i(i_s_23),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_24(.data_o(o_s_24),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_24),.data_i(i_s_24),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_25(.data_o(o_s_25),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_25),.data_i(i_s_25),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_26(.data_o(o_s_26),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_26),.data_i(i_s_26),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_27(.data_o(o_s_27),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_27),.data_i(i_s_27),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_28(.data_o(o_s_28),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_28),.data_i(i_s_28),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_29(.data_o(o_s_29),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_29),.data_i(i_s_29),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_30(.data_o(o_s_30),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_30),.data_i(i_s_30),.oen_i(!wen_1));
tq_ram_1p_16x32  #(.Addr_Width(5), .Word_Width(16)) ram_1p_31(.data_o(o_s_31),.clk(clk),.cen_i(!enable_0),.wen_i(wen_0),.addr_i(add_31),.data_i(i_s_31),.oen_i(!wen_1));

endmodule